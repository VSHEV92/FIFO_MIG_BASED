// ------------------------------------------------------
//-------------------- тестовый набор x2 ----------------
// ------------------------------------------------------
parameter int PHY_to_UI_Rate = 2; // 1 - X4, 2 - X2
parameter int Max_Burst_Len = 16;
parameter int RW_Delay_Value = 4;
parameter int Base_Address = 400;
parameter int Memory_Size = 100;
parameter int MIG_Data_Port_Size = 64;
parameter int MIG_Addr_Port_Size = 28;
parameter int IO_Fifo_Depth = 32;
